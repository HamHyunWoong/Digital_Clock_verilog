module state_mod(input clk, input btn1,output clk_out,output selectout);


reg tap;
reg game_select;

assign

assign selectout = game_select;
assign clk_out = tap;



endmodule